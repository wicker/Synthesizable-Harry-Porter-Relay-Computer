/* Author: Jenner Hanni
 * Project: Harry Porter Relay Computer
 * File: The ALU, which uses eight 1-bit logic blocks which
 * can compute logical AND, OR, XOR, and NOT on all 8 bits.
 * License: MIT http://opensource.org/licenses/MIT
*/

module ALU (input [7:0] b, c, output [7:0] result);

  wire AND, OR, XOR, NOT;
  reg AND_var, OR_var, XOR_var, NOT_var;

  // 
  // 3-to-8 Function Decoder
  // 
 
endmodule
