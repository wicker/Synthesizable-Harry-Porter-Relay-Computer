/* Author: Jenner Hanni
 * Project: Harry Porter Relay Computer
 * File: Result Bus Interface
 * License: MIT http://opensource.org/licenses/MIT
*/

module ResultBus (input logic [7:0] result, output [7:0] alu_result);

  

endmodule
