/* Author: Jenner Hanni
 * Project: Harry Porter Relay Computer
 * File: Register unit
 * License: MIT http://opensource.org/licenses/MIT
*/
