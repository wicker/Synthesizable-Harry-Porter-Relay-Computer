/* Relay testbench */
